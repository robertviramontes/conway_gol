//Legal Notice: (C)2014 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module lt24_qsys_nios2_gen2_0_cpu_oci_test_bench (
                                                   // inputs:
                                                    dct_buffer,
                                                    dct_count,
                                                    test_ending,
                                                    test_has_ended
                                                 )
;

  input   [ 29: 0] dct_buffer;
  input   [  3: 0] dct_count;
  input            test_ending;
  input            test_has_ended;


endmodule

